module seq_multiplier ( 
    input logic [15:0] M,
    input logic [15:0] Q,
    input logic clk,
    input logic reset,
    input logic enable,
    output logic [31:0] acc 


)

endmodule